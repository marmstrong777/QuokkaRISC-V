package QuokkaRvPkg;

    typedef enum logic [1:0] {
        MEM_W_SIZE_WORD,
        MEM_W_SIZE_HALF,
        MEM_W_SIZE_BYTE
    } mem_w_size_e;
endpackage